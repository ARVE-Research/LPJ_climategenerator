netcdf CanESM5 {
dimensions:
	lon = 720 ;
	lat = 360 ;
	time = 12 ;
variables:
	double lon(lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:actual_range = -180., 180. ;
		lon:_Storage = "contiguous" ;
		lon:_Storage = "contiguous" ;
		lon:_Endianness = "little" ;
	double lat(lat) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:actual_range = -90., 90. ;
		lat:_Storage = "contiguous" ;
		lat:_Storage = "contiguous" ;
		lat:_Endianness = "little" ;
	double time(time) ;
		time:climatology = "climatology_bounds" ;
		time:avg_period = "0000-01-00 00:00:00" ;
		time:long_name = "time" ;
		time:actual_range = 0., 0. ;
		time:delta_t = "0000-01-00 00:00:00" ;
		time:standard_name = "time" ;
		time:coordinate_defines = "start" ;
		time:calendar = "standard" ;
		time:note = "time coordinate refers to first day of month" ;
		time:units = "days since 0001-01-01 00:00:00" ;
		time:_Storage = "contiguous" ;
		time:_Endianness = "little" ;
	short elv(lat, lon) ;
		elv:long_name = "Elevation above mean sea level" ;
		elv:units = "m" ;
		elv:scale_factor = 1.f ;
		elv:add_offset = 0.f ;
		elv:_FillValue = -32768s ;
		elv:missing_value = -32768s ;
		elv:source = "WorldClim 1.4" ;
		elv:_ChunkSizes = 360, 720 ;
		elv:_DeflateLevel = 1 ;
		elv:valid_range = -353s, 6241s ;
		elv:_Storage = "chunked" ;
		elv:_ChunkSizes = 360, 720 ;
		elv:_DeflateLevel = 1 ;
		elv:_Endianness = "little" ;
	short tmp(time, lat, lon) ;
		tmp:long_name = "Mean temperature" ;
		tmp:units = "degC" ;
		tmp:scale_factor = 0.1f ;
		tmp:add_offset = 0.f ;
		tmp:missing_value = -32768s ;
		tmp:avg_period = "1979-2013" ;
		tmp:source = "CHELSA 1.2" ;
		tmp:_ChunkSizes = 1, 348, 720 ;
		tmp:_DeflateLevel = 1 ;
		tmp:_Endianness = "little" ;
		tmp:valid_range = -640s, 400s ;
		tmp:_Storage = "chunked" ;
		tmp:_Endianness = "little" ;
	short dtr(time, lat, lon) ;
		dtr:long_name = "Diurnal temperature range" ;
		dtr:units = "degC" ;
		dtr:scale_factor = 0.1f ;
		dtr:add_offset = 0.f ;
		dtr:_FillValue = -32768s ;
		dtr:missing_value = -32768s ;
		dtr:avg_period = "1979-2013" ;
		dtr:source = "CHELSA 1.2" ;
		dtr:_ChunkSizes = 1, 348, 720 ;
		dtr:_DeflateLevel = 1 ;
		dtr:valid_range = -24s, 272s ;
		dtr:_Storage = "chunked" ;
		dtr:_Endianness = "little" ;
	short pre(time, lat, lon) ;
		pre:long_name = "Total precipitation" ;
		pre:units = "mm" ;
		pre:scale_factor = 1.f ;
		pre:add_offset = 0. ;
		pre:missing_value = -32768s ;
		pre:avg_period = "1979-2013" ;
		pre:source = "CHELSA 1.2" ;
		pre:_ChunkSizes = 1, 348, 720 ;
		pre:_DeflateLevel = 1 ;
		pre:valid_range = -32767s, 2500s ;
		pre:_Storage = "chunked" ;
		pre:_Endianness = "little" ;
	short wet(time, lat, lon) ;
		wet:long_name = "Number of days with >0.1 mm precipitation per month" ;
		wet:units = "days" ;
		wet:scale_factor = 0.1f ;
		wet:add_offset = 0.f ;
		wet:_FillValue = -32768s ;
		wet:missing_value = -32768s ;
		wet:avg_period = "1979-2013" ;
		wet:source = "CHELSEA 1.2+" ;
		wet:_ChunkSizes = 1, 348, 720 ;
		wet:_DeflateLevel = 1 ;
		wet:valid_range = 0s, 310s ;
		wet:_Storage = "chunked" ;
		wet:_Endianness = "little" ;
	short cld(time, lat, lon) ;
		cld:long_name = "percent of sky covered by clouds" ;
		cld:units = "percent" ;
		cld:scale_factor = 0.01f ;
		cld:add_offset = 0.f ;
		cld:_FillValue = -32768s ;
		cld:missing_value = -32768s ;
		cld:avg_period = "2000-2014" ;
		cld:source = "MODCF 1-km cloud climatology" ;
		cld:_ChunkSizes = 1, 348, 720 ;
		cld:_DeflateLevel = 1 ;
		cld:valid_range = -353s, 10000s ;
		cld:_Storage = "chunked" ;
		cld:_Endianness = "little" ;
	short wnd(time, lat, lon) ;
		wnd:long_name = "10m windspeed" ;
		wnd:units = "m s-1" ;
		wnd:scale_factor = 0.01f ;
		wnd:add_offset = 0.f ;
		wnd:_FillValue = -32768s ;
		wnd:missing_value = -32768s ;
		wnd:avg_period = "1961-1990" ;
		wnd:source = "CRU CL 2.00" ;
		wnd:_ChunkSizes = 1, 348, 720 ;
		wnd:_DeflateLevel = 1 ;
		wnd:valid_range = 10s, 980s ;
		wnd:_Storage = "chunked" ;
		wnd:_Endianness = "little" ;
	float lght(time, lat, lon) ;
		lght:long_name = "cloud-to-ground lightning strikes" ;
		lght:units = "strikes km-2 d-1" ;
		lght:scale_factor = 1.f ;
		lght:add_offset = 0.f ;
		lght:_FillValue = -32768.f ;
		lght:missing_value = -32768.f ;
		lght:avg_period = "2010-2019" ;
		lght:source = "WLLN monthly lightning flashes" ;
		lght:_ChunkSizes = 1, 348, 720 ;
		lght:_DeflateLevel = 1 ;
		lght:valid_range = 0., 32150.f ;
		lght:_Storage = "chunked" ;
		lght:_Endianness = "little" ;

// global attributes:
		:Conventions = "COARDS, CF-1.0" ;
		:title = "Hybrid long-term mean climatology for global land areas, 30 minute degree grid, v. 1.0" ;
		:note = "30 minute data created by taking median values from 5min WorldClim data and 10min CRU data" ;
		:node_offset = 1 ;
		:history = "Thu Jul  9 22:07:29 2015: ncatted -a units,time,o,c,days since 0001-01-01 00:00:00 climate_wwna_shelves.nc" ;
		:_SuperblockVersion = 2 ;
		:_IsNetcdf4 = 1 ;
		:_Format = "netCDF-4" ;
data:

 lon = -179.75, -179.25, -178.75, -178.25, -177.75, -177.25, -176.75, 
    -176.25, -175.75, -175.25, -174.75, -174.25, -173.75, -173.25, -172.75, 
    -172.25, -171.75, -171.25, -170.75, -170.25, -169.75, -169.25, -168.75, 
    -168.25, -167.75, -167.25, -166.75, -166.25, -165.75, -165.25, -164.75, 
    -164.25, -163.75, -163.25, -162.75, -162.25, -161.75, -161.25, -160.75, 
    -160.25, -159.75, -159.25, -158.75, -158.25, -157.75, -157.25, -156.75, 
    -156.25, -155.75, -155.25, -154.75, -154.25, -153.75, -153.25, -152.75, 
    -152.25, -151.75, -151.25, -150.75, -150.25, -149.75, -149.25, -148.75, 
    -148.25, -147.75, -147.25, -146.75, -146.25, -145.75, -145.25, -144.75, 
    -144.25, -143.75, -143.25, -142.75, -142.25, -141.75, -141.25, -140.75, 
    -140.25, -139.75, -139.25, -138.75, -138.25, -137.75, -137.25, -136.75, 
    -136.25, -135.75, -135.25, -134.75, -134.25, -133.75, -133.25, -132.75, 
    -132.25, -131.75, -131.25, -130.75, -130.25, -129.75, -129.25, -128.75, 
    -128.25, -127.75, -127.25, -126.75, -126.25, -125.75, -125.25, -124.75, 
    -124.25, -123.75, -123.25, -122.75, -122.25, -121.75, -121.25, -120.75, 
    -120.25, -119.75, -119.25, -118.75, -118.25, -117.75, -117.25, -116.75, 
    -116.25, -115.75, -115.25, -114.75, -114.25, -113.75, -113.25, -112.75, 
    -112.25, -111.75, -111.25, -110.75, -110.25, -109.75, -109.25, -108.75, 
    -108.25, -107.75, -107.25, -106.75, -106.25, -105.75, -105.25, -104.75, 
    -104.25, -103.75, -103.25, -102.75, -102.25, -101.75, -101.25, -100.75, 
    -100.25, -99.75, -99.25, -98.75, -98.25, -97.75, -97.25, -96.75, -96.25, 
    -95.75, -95.25, -94.75, -94.25, -93.75, -93.25, -92.75, -92.25, -91.75, 
    -91.25, -90.75, -90.25, -89.75, -89.25, -88.75, -88.25, -87.75, -87.25, 
    -86.75, -86.25, -85.75, -85.25, -84.75, -84.25, -83.75, -83.25, -82.75, 
    -82.25, -81.75, -81.25, -80.75, -80.25, -79.75, -79.25, -78.75, -78.25, 
    -77.75, -77.25, -76.75, -76.25, -75.75, -75.25, -74.75, -74.25, -73.75, 
    -73.25, -72.75, -72.25, -71.75, -71.25, -70.75, -70.25, -69.75, -69.25, 
    -68.75, -68.25, -67.75, -67.25, -66.75, -66.25, -65.75, -65.25, -64.75, 
    -64.25, -63.75, -63.25, -62.75, -62.25, -61.75, -61.25, -60.75, -60.25, 
    -59.75, -59.25, -58.75, -58.25, -57.75, -57.25, -56.75, -56.25, -55.75, 
    -55.25, -54.75, -54.25, -53.75, -53.25, -52.75, -52.25, -51.75, -51.25, 
    -50.75, -50.25, -49.75, -49.25, -48.75, -48.25, -47.75, -47.25, -46.75, 
    -46.25, -45.75, -45.25, -44.75, -44.25, -43.75, -43.25, -42.75, -42.25, 
    -41.75, -41.25, -40.75, -40.25, -39.75, -39.25, -38.75, -38.25, -37.75, 
    -37.25, -36.75, -36.25, -35.75, -35.25, -34.75, -34.25, -33.75, -33.25, 
    -32.75, -32.25, -31.75, -31.25, -30.75, -30.25, -29.75, -29.25, -28.75, 
    -28.25, -27.75, -27.25, -26.75, -26.25, -25.75, -25.25, -24.75, -24.25, 
    -23.75, -23.25, -22.75, -22.25, -21.75, -21.25, -20.75, -20.25, -19.75, 
    -19.25, -18.75, -18.25, -17.75, -17.25, -16.75, -16.25, -15.75, -15.25, 
    -14.75, -14.25, -13.75, -13.25, -12.75, -12.25, -11.75, -11.25, -10.75, 
    -10.25, -9.75, -9.25, -8.75, -8.25, -7.75, -7.25, -6.75, -6.25, -5.75, 
    -5.25, -4.75, -4.25, -3.75, -3.25, -2.75, -2.25, -1.75, -1.25, -0.75, 
    -0.25, 0.25, 0.75, 1.25, 1.75, 2.25, 2.75, 3.25, 3.75, 4.25, 4.75, 5.25, 
    5.75, 6.25, 6.75, 7.25, 7.75, 8.25, 8.75, 9.25, 9.75, 10.25, 10.75, 
    11.25, 11.75, 12.25, 12.75, 13.25, 13.75, 14.25, 14.75, 15.25, 15.75, 
    16.25, 16.75, 17.25, 17.75, 18.25, 18.75, 19.25, 19.75, 20.25, 20.75, 
    21.25, 21.75, 22.25, 22.75, 23.25, 23.75, 24.25, 24.75, 25.25, 25.75, 
    26.25, 26.75, 27.25, 27.75, 28.25, 28.75, 29.25, 29.75, 30.25, 30.75, 
    31.25, 31.75, 32.25, 32.75, 33.25, 33.75, 34.25, 34.75, 35.25, 35.75, 
    36.25, 36.75, 37.25, 37.75, 38.25, 38.75, 39.25, 39.75, 40.25, 40.75, 
    41.25, 41.75, 42.25, 42.75, 43.25, 43.75, 44.25, 44.75, 45.25, 45.75, 
    46.25, 46.75, 47.25, 47.75, 48.25, 48.75, 49.25, 49.75, 50.25, 50.75, 
    51.25, 51.75, 52.25, 52.75, 53.25, 53.75, 54.25, 54.75, 55.25, 55.75, 
    56.25, 56.75, 57.25, 57.75, 58.25, 58.75, 59.25, 59.75, 60.25, 60.75, 
    61.25, 61.75, 62.25, 62.75, 63.25, 63.75, 64.25, 64.75, 65.25, 65.75, 
    66.25, 66.75, 67.25, 67.75, 68.25, 68.75, 69.25, 69.75, 70.25, 70.75, 
    71.25, 71.75, 72.25, 72.75, 73.25, 73.75, 74.25, 74.75, 75.25, 75.75, 
    76.25, 76.75, 77.25, 77.75, 78.25, 78.75, 79.25, 79.75, 80.25, 80.75, 
    81.25, 81.75, 82.25, 82.75, 83.25, 83.75, 84.25, 84.75, 85.25, 85.75, 
    86.25, 86.75, 87.25, 87.75, 88.25, 88.75, 89.25, 89.75, 90.25, 90.75, 
    91.25, 91.75, 92.25, 92.75, 93.25, 93.75, 94.25, 94.75, 95.25, 95.75, 
    96.25, 96.75, 97.25, 97.75, 98.25, 98.75, 99.25, 99.75, 100.25, 100.75, 
    101.25, 101.75, 102.25, 102.75, 103.25, 103.75, 104.25, 104.75, 105.25, 
    105.75, 106.25, 106.75, 107.25, 107.75, 108.25, 108.75, 109.25, 109.75, 
    110.25, 110.75, 111.25, 111.75, 112.25, 112.75, 113.25, 113.75, 114.25, 
    114.75, 115.25, 115.75, 116.25, 116.75, 117.25, 117.75, 118.25, 118.75, 
    119.25, 119.75, 120.25, 120.75, 121.25, 121.75, 122.25, 122.75, 123.25, 
    123.75, 124.25, 124.75, 125.25, 125.75, 126.25, 126.75, 127.25, 127.75, 
    128.25, 128.75, 129.25, 129.75, 130.25, 130.75, 131.25, 131.75, 132.25, 
    132.75, 133.25, 133.75, 134.25, 134.75, 135.25, 135.75, 136.25, 136.75, 
    137.25, 137.75, 138.25, 138.75, 139.25, 139.75, 140.25, 140.75, 141.25, 
    141.75, 142.25, 142.75, 143.25, 143.75, 144.25, 144.75, 145.25, 145.75, 
    146.25, 146.75, 147.25, 147.75, 148.25, 148.75, 149.25, 149.75, 150.25, 
    150.75, 151.25, 151.75, 152.25, 152.75, 153.25, 153.75, 154.25, 154.75, 
    155.25, 155.75, 156.25, 156.75, 157.25, 157.75, 158.25, 158.75, 159.25, 
    159.75, 160.25, 160.75, 161.25, 161.75, 162.25, 162.75, 163.25, 163.75, 
    164.25, 164.75, 165.25, 165.75, 166.25, 166.75, 167.25, 167.75, 168.25, 
    168.75, 169.25, 169.75, 170.25, 170.75, 171.25, 171.75, 172.25, 172.75, 
    173.25, 173.75, 174.25, 174.75, 175.25, 175.75, 176.25, 176.75, 177.25, 
    177.75, 178.25, 178.75, 179.25, 179.75 ;

 lat = -89.75, -89.25, -88.75, -88.25, -87.75, -87.25, -86.75, -86.25, 
    -85.75, -85.25, -84.75, -84.25, -83.75, -83.25, -82.75, -82.25, -81.75, 
    -81.25, -80.75, -80.25, -79.75, -79.25, -78.75, -78.25, -77.75, -77.25, 
    -76.75, -76.25, -75.75, -75.25, -74.75, -74.25, -73.75, -73.25, -72.75, 
    -72.25, -71.75, -71.25, -70.75, -70.25, -69.75, -69.25, -68.75, -68.25, 
    -67.75, -67.25, -66.75, -66.25, -65.75, -65.25, -64.75, -64.25, -63.75, 
    -63.25, -62.75, -62.25, -61.75, -61.25, -60.75, -60.25, -59.75, -59.25, 
    -58.75, -58.25, -57.75, -57.25, -56.75, -56.25, -55.75, -55.25, -54.75, 
    -54.25, -53.75, -53.25, -52.75, -52.25, -51.75, -51.25, -50.75, -50.25, 
    -49.75, -49.25, -48.75, -48.25, -47.75, -47.25, -46.75, -46.25, -45.75, 
    -45.25, -44.75, -44.25, -43.75, -43.25, -42.75, -42.25, -41.75, -41.25, 
    -40.75, -40.25, -39.75, -39.25, -38.75, -38.25, -37.75, -37.25, -36.75, 
    -36.25, -35.75, -35.25, -34.75, -34.25, -33.75, -33.25, -32.75, -32.25, 
    -31.75, -31.25, -30.75, -30.25, -29.75, -29.25, -28.75, -28.25, -27.75, 
    -27.25, -26.75, -26.25, -25.75, -25.25, -24.75, -24.25, -23.75, -23.25, 
    -22.75, -22.25, -21.75, -21.25, -20.75, -20.25, -19.75, -19.25, -18.75, 
    -18.25, -17.75, -17.25, -16.75, -16.25, -15.75, -15.25, -14.75, -14.25, 
    -13.75, -13.25, -12.75, -12.25, -11.75, -11.25, -10.75, -10.25, -9.75, 
    -9.25, -8.75, -8.25, -7.75, -7.25, -6.75, -6.25, -5.75, -5.25, -4.75, 
    -4.25, -3.75, -3.25, -2.75, -2.25, -1.75, -1.25, -0.75, -0.25, 0.25, 
    0.75, 1.25, 1.75, 2.25, 2.75, 3.25, 3.75, 4.25, 4.75, 5.25, 5.75, 6.25, 
    6.75, 7.25, 7.75, 8.25, 8.75, 9.25, 9.75, 10.25, 10.75, 11.25, 11.75, 
    12.25, 12.75, 13.25, 13.75, 14.25, 14.75, 15.25, 15.75, 16.25, 16.75, 
    17.25, 17.75, 18.25, 18.75, 19.25, 19.75, 20.25, 20.75, 21.25, 21.75, 
    22.25, 22.75, 23.25, 23.75, 24.25, 24.75, 25.25, 25.75, 26.25, 26.75, 
    27.25, 27.75, 28.25, 28.75, 29.25, 29.75, 30.25, 30.75, 31.25, 31.75, 
    32.25, 32.75, 33.25, 33.75, 34.25, 34.75, 35.25, 35.75, 36.25, 36.75, 
    37.25, 37.75, 38.25, 38.75, 39.25, 39.75, 40.25, 40.75, 41.25, 41.75, 
    42.25, 42.75, 43.25, 43.75, 44.25, 44.75, 45.25, 45.75, 46.25, 46.75, 
    47.25, 47.75, 48.25, 48.75, 49.25, 49.75, 50.25, 50.75, 51.25, 51.75, 
    52.25, 52.75, 53.25, 53.75, 54.25, 54.75, 55.25, 55.75, 56.25, 56.75, 
    57.25, 57.75, 58.25, 58.75, 59.25, 59.75, 60.25, 60.75, 61.25, 61.75, 
    62.25, 62.75, 63.25, 63.75, 64.25, 64.75, 65.25, 65.75, 66.25, 66.75, 
    67.25, 67.75, 68.25, 68.75, 69.25, 69.75, 70.25, 70.75, 71.25, 71.75, 
    72.25, 72.75, 73.25, 73.75, 74.25, 74.75, 75.25, 75.75, 76.25, 76.75, 
    77.25, 77.75, 78.25, 78.75, 79.25, 79.75, 80.25, 80.75, 81.25, 81.75, 
    82.25, 82.75, 83.25, 83.75, 84.25, 84.75, 85.25, 85.75, 86.25, 86.75, 
    87.25, 87.75, 88.25, 88.75, 89.25, 89.75 ;

 time = 0, 31, 59, 90, 120, 151, 181, 212, 243, 273, 304, 334 ;
}
